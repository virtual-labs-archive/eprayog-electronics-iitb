Full Wave Rectifier

.MODEL DIO D( IS=1.8E-14 RS=2 BV=50.0 IBV=1e-4
+ CJO=2e-12  M=0.333 N=2.06 TT=4.32e-9)

Rs 1 2 .5
Lp 2 0 1mH
Ls1 3 0 1mH
Ls2 0 4 1mH
D1 3 5 DIO
D2 4 5 DIO
R2 5 0 5K
Kps  Lp  Ls1  1
Kps1  Lp  Ls2  1
Kss  Ls1  Ls2  1

C1 5 0 5u

v1 1 0 sin(0 25V 1k)

.tran 0.01m 5m

.control

run
plot v(1) v(5)

.endc

.end
