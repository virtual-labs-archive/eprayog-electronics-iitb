**bjt inverter
.model bjt npn (is=10e-16, bf=220, va=50v, cje=20p, cjc=25p)
V1 1 0 dc 10
Rb 1 2 20k
Rc 4 3 12k
Q1 3 2 0 BJT
V2 4 0 dc 5
.dc v1 0 5 0.5
.control
run
plot v(3) v(1)

.endc
.end
