DIODE I-V CURVE AT T=300K
.MODEL DIO D( IS=1.8E-10 RS=2 BV=50.0 IBV=1e-4+ CJO=1e-12 M=0.333 N=2.06 TT=4.32e-9 VJ=1e-6)
.TEMP 27

D1 3 0 DIO
R1 1 2 100
V1 1 0 dc 0v
Vmeas 2 3 dc 0
.dc v1 0 5 0.2

.control
run
plot i(vmeas) vs v(3)
.endc
.end
